// 2024.9.23 Epi Week 2 code 6
// target: simulate WIRE
module top_module(input in, output out);
    assign out = in;
endmodule