// 2024.9.23 Epi Week 2 code 1
// target: No input, output 0

module top_module(output zero);
    assign zero = 0;
endmodule