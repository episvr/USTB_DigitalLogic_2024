// 2024.9.23 Epi Week 2 code 2
// target: NOT gate
module top_module(input in, output out);
    assign out = ~in;
endmodule